import uvm_pkg::*;
import riscv_txn_pkg::*;
import pc_tb_pkg::*;

`include "uvm_macros.svh"

class rf_test extends uvm_test;

  `uvm_component_utils(rf_test)

  rf_env env;

  function new(string name = "rf_test", uvm_component parent);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = rf_env::type_id::create("env", this);
  endfunction

  virtual task run_phase(uvm_phase phase);

    rf_base_sequence seq;

    phase.raise_objection(this);

    seq = rf_base_sequence::type_id::create("seq");

    seq.start(env.agent.sequencer);

    phase.drop_objection(this);

  endtask

endclass