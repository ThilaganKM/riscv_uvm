import uvm_pkg::*;
`include "uvm_macros.svh"
module tb_top;

    //--------------------------------------------------
    // Clock
    //--------------------------------------------------

    logic clk;

    always #5 clk = ~clk;

    //--------------------------------------------------
    // Interface
    //--------------------------------------------------

    pc_if pcif(clk);

    //--------------------------------------------------
    // DUT
    //--------------------------------------------------

    pc dut (
        .clk    (clk),
        .reset  (pcif.reset),
        .en     (pcif.en),
        .PCNext (pcif.PCNext),
        .PC     (pcif.PC)
    );

    //--------------------------------------------------
    // UVM Configuration
    //--------------------------------------------------

    initial begin

        //--------------------------------------------------
        // Initialize Clock
        //--------------------------------------------------

        clk = 0;

        //--------------------------------------------------
        // Pass Interface to UVM
        //--------------------------------------------------

        uvm_config_db #(virtual pc_if)::set(
            null,
            "*",
            "vif",
            pcif
        );

        //--------------------------------------------------
        // Run Test
        //--------------------------------------------------

        run_test("pc_test");

    end

endmodule