package pipeline_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "pipeline_scoreboard.sv"
  `include "riscv_rand_instr.sv"
  `include "pipeline_env.sv"
  `include "pipeline_test.sv"

endpackage