class fwd_sequencer extends uvm_sequencer #(fwd_seq_item);

  `uvm_component_utils(fwd_sequencer)

  function new(string name = "fwd_sequencer", uvm_component parent);
    super.new(name, parent);
  endfunction

endclass