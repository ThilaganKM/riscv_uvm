class data_mem_sequencer extends uvm_sequencer #(dmem_seq_item);
  `uvm_component_utils(data_mem_sequencer)
  function new(string name, uvm_component parent);
    super.new(name,parent);
  endfunction
endclass