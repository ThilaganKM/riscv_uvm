class control_unit_env extends uvm_env;

  `uvm_component_utils(control_unit_env)

  control_unit_agent      agent;
  control_unit_scoreboard sb;

  function new(string name = "control_unit_env", uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    agent = control_unit_agent::type_id::create("agent", this);
    sb    = control_unit_scoreboard::type_id::create("sb", this);

  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);

    agent.mon.ap.connect(sb.analysis_export);

  endfunction

endclass